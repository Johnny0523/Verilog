module Test2(clk,enable,seed,D);

input clk,enable,seed;
output [5:0]D;

reg [5:0]D;

always @(posedge clk)
begin
	if(enable)
	begin
	D[0]<=seed;
	D[1]<=D[0];
	D[2]<=D[1];
	D[3]<=D[2];
	D[4]<=D[3];
	D[5]<=D[4];
	end
	else
	begin;
	D[0]<=D[4]^D[5];
	D[1]<=D[0];
	D[2]<=D[1];
	D[3]<=D[2];
	D[4]<=D[3];
	D[5]<=D[4];
	end
end
endmodule